int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
int sum(int a, int b) {
	int c = a+b;
	return c;
}

void main() {
	int x = 5;
	int y = 10;
	
	int c = sum(x, y);
	
	if(c > 50) {
		c = c + 1;
	}
}
