void main() {
	int x = 5;
	int y = 10;

	int z = x + y;
}