void main() {
	Array[Array[int, 3], 3] a = [[0, 1, 2], [3, 4, 5], [6, 7, 8]];
}